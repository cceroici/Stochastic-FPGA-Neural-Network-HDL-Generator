


module NN_GRADCALC(delta,a,dalpha);

input delta,a;

output dalpha;

and a0(dalpha,delta,a);

endmodule